module dev_in(data_in, data_out);
  input [31:0] data_in;
  output [31:0] data_out;
  
  assign data_out = data_in;
  
endmodule
